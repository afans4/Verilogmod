module multde (
    input clk,
    input [7:0] data,
    input rstn,
    output [7:0] odata
);
    parameter K = 13'b0_01_0010_1000_11;
endmodule //multde