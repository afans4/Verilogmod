`timescale 1ps/1ps
//  Module: text

module tb_jiajian;
    reg        [2:0] a,b,c;
    reg signed [2:0] sa,sb,sc;
    reg        [3:0] sum;
    reg signed [3:0] ssum;
    reg        [2:0] us;
    reg signed [2:0] ss;
    initial begin
        a = 3'b110;
        b = 3'b010;
        c = 3'b111;
        sa = 3'b110;
        sb = 3'b010;
        sc = 3'b111;
        $display("-----------------------");
        $display("-");
        $display("ssum is signed");
        ssum = sb-sa;
        $display("1:S%b - S%b = %b", sb,sa,ssum);
        ssum = sb - a;
        $display("2:S%b - %b = %b", sb,a,ssum);
        ssum = sb-sa;
        $display("3:S%b -S%b = %b", sb,sa,ssum);
        ssum = b-sa;
        $display("4:%b - S%b = %b", b,sa,ssum);
        $display("-----------------------");
        $display("sum is unsigned");
        sum = sb-sa;
        $display("1:S%b - S%b = %b", sb,sa,sum);
        sum = sb - a;
        $display("2:S%b - %b = %b", sb,a,sum);
        sum = sb-sa;
        $display("3:S%b - S%b = %b", sb,sa,sum);
        sum = b-sa;
        $display("4:%b - S%b = %b", b,sa,sum);
        $display("-----------------------");
        $display("+");
        $display("ssum is signed");
        ssum = sb+sc;
        $display("1:S%b + S%b = %b", sb,sc,ssum);
        ssum = sb + c;
        $display("2:S%b + %b = %b", sb,c,ssum);
        ssum = sb+sc;
        $display("3:S%b +S%b = %b", sb,sc,ssum);
        ssum = b+sc;
        $display("4:%b + S%b = %b", b,sc,ssum);
        $display("-----------------------");
        $display("sum is unsigned");
        sum = sb+sc;
        $display("1:S%b + S%b = %b", sb,sc,sum);
        sum = sb + c;
        $display("2:S%b + %b = %b", sb,c,sum);
        sum = sb+sc;
        $display("3:S%b + S%b = %b", sb,sc,sum);
        sum = b+sc;
        $display("4:%b + S%b = %b", b,sc,sum);
        $display("-----------------------");
        a = 3'b001;
        b = 3'b100;
        sum = a-b;
        us = a-b;
        ss = a-b;
        $display("%b - %b = %b",a,b,sum);
        $display("us = %b,ss = %b",us,ss);
        $display("--------------------------");
        a = 3'b101;
        sa = 3'b101;
        b = 3'b011;
        sb = 3'b011;
        c = a >>> 1;
        sc = a >>> 1;
        $display("%0b >>> 1 = s%b",a,sc);
        $display("%0b >>> 1 = %b",a,c);
        $display("--------------------------");
        c = sa >>> 1;
        sc = sa >>> 1;
        $display("s%b >>> 1 = s%b",sa,sc);
        $display("s%b >>> 1 = %b",sa,c);
        $display("--------------------------");
        c = b >>> 1;
        sc = b >>> 1;
        $display("%b >>> 1 = s%b",b,sc);
        $display("%b >>> 1 = %b",b,c);
        $display("--------------------------");
        c = sb >>> 1;
        sc = sb >>> 1;
        $display("s%b >>> 1 = s%b",sb,sc);
        $display("s%b >>> 1 = %b",sb,c);
        $display("--------------------------");
        $stop();
    end
    
endmodule
