//-----------------------------------------------------------------
//Copyright (c) 2014-2020 All rights reserved
//Author  : 383423151@qq.com
//File    : center512
//Create  : 2021-07-21
//Revise  : 2021-
//Editor  : Vscode,tab size (4)
//Funciton:
//
//------------------------------------------------------------------
module center512(
    input clk,
    input rstn,
    input [7:0] idata,
    input en_in,
    output [7:0] max_data,
    output [8:0] max_id,
    output [8:0] cent_id,
    output en_out
    );

    
endmodule: center512
