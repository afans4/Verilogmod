`include "uvm_macros.svh"
import uvm_pkg::*;

`include "dut_if.sv"
`include "transaction_i.sv"
`include "transaction_o.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "remodel.sv"
`include "scoreboard.sv"
`include "my_env.sv"
`include "base_test.sv"
`include "my_case0.sv"
