class myclass;
    bit [7:0] data;
    string name;
    function new(string name);
        this.name = name;
    endfunction
endclass
