module fifo (
    input clk,
    input rstn,
    input 
);

endmodule //fifo